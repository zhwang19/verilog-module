library verilog;
use verilog.vl_types.all;
entity tb_pipeline_mul is
end tb_pipeline_mul;
