library verilog;
use verilog.vl_types.all;
entity tb_synch_fifo is
end tb_synch_fifo;
