library verilog;
use verilog.vl_types.all;
entity tb_tb_binary_to_gray is
end tb_tb_binary_to_gray;
