library verilog;
use verilog.vl_types.all;
entity tb_clk_float_divider is
end tb_clk_float_divider;
