library verilog;
use verilog.vl_types.all;
entity tb_divider is
end tb_divider;
