library verilog;
use verilog.vl_types.all;
entity tb_sequence_mul is
end tb_sequence_mul;
