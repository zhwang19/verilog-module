library verilog;
use verilog.vl_types.all;
entity tb_avoid_fluttering is
end tb_avoid_fluttering;
