library verilog;
use verilog.vl_types.all;
entity tb_spi_module is
end tb_spi_module;
