library verilog;
use verilog.vl_types.all;
entity tb_uart_top is
end tb_uart_top;
