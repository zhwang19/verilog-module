library verilog;
use verilog.vl_types.all;
entity tb_syn_shaping is
end tb_syn_shaping;
