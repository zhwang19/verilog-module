library verilog;
use verilog.vl_types.all;
entity tb_gray_to_binary is
end tb_gray_to_binary;
